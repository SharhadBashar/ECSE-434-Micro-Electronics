Experiment 1.2
*Circuit description*

*Power sources*
Vin 0 1 AC 1m 0
Vcc 6 0 DC 5
Vee 7 0 DC -5

*Elements*
C1 1 2 1uF
R1 2 0 150K
Rpot 4 0 5K
R2 5 4 750K
X1 2 4 6 7 5 TL084

**ANALYSIS REQUUEST**
.AC DEC 3 0.1Hz 1MegHz

**OUTPUT REQUEST**
*.PLOT TRAN V(6) V(1)
.PROBE 


**TL084**
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt TL084    1 2 3 4 5
*
x_tl084 1 2 3 4 5 TL082
.ends




**TL082**
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt TL082    1 2 3 4 5
*
c1   11 12 2.412E-12
c2    6  7 18.00E-12
css  10 99 5.400E-12
dc    5 53 dy
de   54  5 dy
dlp  90 91 dx
dln  92 90 dx
dp    4  3 dx
egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
fb    7 99 poly(5) vb vc ve vlp vln 0 3.467E6 -1E3 1E3 3E6 -3E6
ga    6  0 11 12 339.3E-6
gcm   0  6 10 99 17.01E-9
iss  10  4 dc 234.0E-6
hlim 90  0 vlim 1K
j1   11  2 10 jx
j2   12  1 10 jx
r2    6  9 100.0E3
rd1   3 11 2.947E3
rd2   3 12 2.947E3
ro1   8  5 50
ro2   7 99 170
rp    3  4 20.00E3
rss  10 99 854.7E3
vb    9  0 dc 0
vc    3 53 dc 1.500
ve   54  4 dc 1.500
vlim  7  8 dc 0
vlp  91  0 dc 50
vln   0 92 dc 50
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx NJF(Is=2.500E-12 Beta=984.2E-6 Vto=-1)
.ends




.END