Prelab 3.1
*Class A Output Stage*

*Sources
Vin 0 1 SIN (0 0.2 10K 0 0 0)
VCC1 4 0 5
VCC2 5 0 5
VEE 3 0 -5

*Elements
*Capacitors
C4 1 2 22u
CL 3 0 22u
CP 4 0 22u
C5 7 8 22u

*Resistors
R10 2 4 4.3K
R11 2 3 5.7K
R12 6 5 48
RL 8 0 8
RE1 3 9 47
RE2 3 10 47 

*Transisors 
QT5 6 6 9 MPS3704
QT6 7 6 10 MPS3704
QT7 4 2 7 MPS3704

.model MPS3704	NPN(Is=26.03f Xti=3 Eg=1.11 Vaf=90.7 Bf=736.1K Ne=1.232
+		Ise=26.03f Ikf=.1983 Xtb=1.5 Br=1.024 Nc=2 Isc=0 Ikr=0 Rc=.5
+		Cjc=11.01p Mjc=.3763 Vjc=.75 Fc=.5 Cje=24.07p Mje=.3641 Vje=.75
+		Tr=233.8n Tf=1.03n Itf=0 Vtf=0 Xtf=0 Rb=10)
*		Motorola	pid=2N4400	case=TO92
*		88-09-13 bam	creation

*Analysis Request
.probe
.TRAN 0.1m 2m

.END