Exp 5.1
**Circuit Description
*Voltage Supply
Vin1 30 0  SIN (0 0.5m 10K)
Vin2 31 0  SIN (0 1 464K)
*Vin 0 30 AC 1m 0
*Vin2 0 31 AC 1m 0

E1_mult 0 2 value {V(30)*V(31)}

XPreamp 2 3 Preamp
XDemod 3 4 Demod
XBBAmp 4 5 BBAmp
XCAOS 5 6 CAOS

*Analysis Request
.PROBE
.TRAN 0 5m
*.AC DEC 10 0.01Hz 10MegHz

*********************** Preamplifier ***************************
.SUBCKT Preamp 1 10
	*Voltage Sources
	*Vin 0 1 AC 1m 0

	VCC 3 0 5V

	*Elements*
	*Capacitors 
	C2 1 2 1u
	C3 3 0 1u
	CB 4 0 1u

	*Resisors
	R5 2 0 22k
	R4 2 3 28k
	R6 3 4 25k
	R7 4 0 70k
	RE 6 0 40
	R9 10 0 100

	*Transisors
	QT1 5 2 6 MPS3704
	QT2 8 4 5 MPS3704
	QT3 3 8 9 MPS3704
	QT4 3 9 10 MPS3704

	.model MPS3704	NPN(Is=26.03f Xti=3 Eg=1.11 Vaf=90.7 Bf=736.1K Ne=1.232
	+		Ise=26.03f Ikf=.1983 Xtb=1.5 Br=1.024 Nc=2 Isc=0 Ikr=0 Rc=.5
	+		Cjc=11.01p Mjc=.3763 Vjc=.75 Fc=.5 Cje=24.07p Mje=.3641 Vje=.75
	+		Tr=233.8n Tf=1.03n Itf=0 Vtf=0 Xtf=0 Rb=10)
	*		Motorola	pid=2N4400	case=TO92
	*		88-09-13 bam	creation

	*TANK
	RL 3 7 10
	LT 7 8 100uH
	CT 3 8 1nF

	*Analysis Request
	*.probe
	*.TRAN 0.1m 0.5m
	*.AC DEC 3 0.1Hz 1000MEGHz
.ENDS Preamp
******************************************************************

************************* Demodulator ****************************
.SUBCKT Demod 2 3
*
	*Circuit Analysis
	*Vin1 0 1 SIN (0 10 10K 0 0 0)
	*Vin2 1 2 SIN (0 25 0.25Meg 0 0 0)

	D 2 3 1N34A

	.MODEL 1N34A D ( bv=75 cjo=0.5e-12 eg=0.67 ibv=18e-3 is=2e-7 rs=7 n=1.3 vj=0.1 m=0.27 )
	Rdem 3 0 200k
	Cdem 3 0 0.934n

	*analysis request
	*.PROBE
	*.TRAN 0 1m
.ENDS Demod
******************************************************************

************************ BaseBand Amp ****************************
.SUBCKT BBAmp 1 4

	*Circuit description*

	*Power sources*
	*Vin 0 1 AC 1m 0
	Vcc 5 0 DC 5
	Vee 6 0 DC -5

	*Elements*
	C1 1 2 1uF
	R1 2 0 150K
	Rpot 0 3 10K
	R2 3 4 50K
	X1 2 3 5 6 4 TL084

	**ANALYSIS REQUUEST**
	*.AC DEC 10 0.01Hz 10MegHz

	**OUTPUT REQUEST**

	*.PROBE 
.ENDS BBAmp
*-----------------------------------------------------------------------------
	**TL084**
	* connections:   non-inverting input
	*                | inverting input
	*                | | positive power supply
	*                | | | negative power supply
	*                | | | | output
	*                | | | | |
	.subckt TL084    1 2 3 4 5
		*
		X_tl084 1 2 3 4 5 TL082
 	.ends

	**TL082**
*-----------------------------------------------------------------------------
	* connections:non-inverting input
	*             | inverting input
	*             | | positive power supply
	*             | | | negative power supply
	*             | | | | output
	*             | | | | |
	.subckt TL082 1 2 3 4 5
		*
		c1   11 12 2.412E-12
		c2    6  7 18.00E-12
		css  10 99 5.400E-12
		dc    5 53 dy
		de   54  5 dy
		dlp  90 91 dx
		dln  92 90 dx
		dp    4  3 dx
		egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
		fb    7 99 poly(5) vb vc ve vlp vln 0 3.467E6 -1E3 1E3 3E6 -3E6
		ga    6  0 11 12 339.3E-6
		gcm   0  6 10 99 17.01E-9
		iss  10  4 dc 234.0E-6
		hlim 90  0 vlim 1K
		j1   11  2 10 jx
		j2   12  1 10 jx
		r2    6  9 100.0E3
		rd1   3 11 2.947E3
		rd2   3 12 2.947E3
		ro1   8  5 50
		ro2   7 99 170
		rp    3  4 20.00E3
		rss  10 99 854.7E3
		vb    9  0 dc 0
		vc    3 53 dc 1.500
		ve   54  4 dc 1.500
		vlim  7  8 dc 0
		vlp  91  0 dc 50
		vln   0 92 dc 50
		.model dx D(Is=800.0E-18 Rs=1)
		.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
		.model jx NJF(Is=2.500E-12 Beta=984.2E-6 Vto=-1)
	.ends
******************************************************************

******************** Class A Output Stage ************************
.SUBCKT CAOS 1 8
	*Class A Output Stage*

	*Sources
	*Vin 0 1 SIN (0 0.2 10K 0 0 0)
	VCC1 4 0 5
	VCC2 5 0 5
	VEE 3 0 -5

	*Elements
	*Capacitors
	C4 1 2 22u
	CL 3 0 22u
	CP 4 0 22u
	C5 7 8 22u

	*Resistors
	R10 2 4 4.3K
	R11 2 3 5.7K
	R12 6 5 48
	RL 8 0 8
	RE1 3 9 47
	RE2 3 10 47 

	*Transisors 
	QT5 6 6 9 MPS3704
	QT6 7 6 10 MPS3704
	QT7 4 2 7 MPS3704

	.model MPS3704	NPN(Is=26.03f Xti=3 Eg=1.11 Vaf=90.7 Bf=736.1K Ne=1.232
	+		Ise=26.03f Ikf=.1983 Xtb=1.5 Br=1.024 Nc=2 Isc=0 Ikr=0 Rc=.5
	+		Cjc=11.01p Mjc=.3763 Vjc=.75 Fc=.5 Cje=24.07p Mje=.3641 Vje=.75
	+		Tr=233.8n Tf=1.03n Itf=0 Vtf=0 Xtf=0 Rb=10)
	*		Motorola	pid=2N4400	case=TO92
	*		88-09-13 bam	creation

	*Analysis Request
	*.probe
	*.TRAN 0.1m 2m

.ENDS CAOS

******************************************************************


.END